module InstructionMemory_P(Address, Instruction);
input [31:0] Address;
output [31:0] Instruction;
reg [31:0] Instruction;
always @(*)
	case(Address[9:2])
		0: Instruction<=32'b00001000000000000000000000000011;	//j Main
		1: Instruction<=32'b00001000000000000000000000100010;	//j Interrupt
		2: Instruction<=32'b000010;	//j Abnormal
		3: Instruction<=32'b00111100000111100100000000000000;	//Main:   lui $fp,16384
		4: Instruction<=32'b00100000000111010000010000000000;	//addi $sp,$zero,1024
		5: Instruction<=32'b10101111110000000000000000001000;	//sw $zero,2($fp)
		6: Instruction<=32'b00100000000010001111100000000000;	//addi $t0,$zero,-2048
		7: Instruction<=32'b10101111110010000000000000000000;	//sw $t0,0($fp)
		8: Instruction<=32'b00100000000010001111111111111111;	//addi $t0,$zero,-1
		9: Instruction<=32'b10101111110010000000000000000100;	//sw $t0,1($fp)
		10:Instruction<=32'b00100000000010000000000000000011;	//addi $t0,$zero,3
		11:Instruction<=32'b10101111110010000000000000001000;	//sw $t0,2($fp)
		12:Instruction<=32'b10001111110010000000000000100000;	//Read1:   lw $t0,8($fp)
		13:Instruction<=32'b00110001000010000000000000001000;	//andi $t0,$t0,8
		14:Instruction<=32'b00010000000010001111111111111101;	//beq $t0,$zero,Read1
		15:Instruction<=32'b10001111110100000000000000011100;	//lw $s0,7($fp)
		16:Instruction<=32'b00000010000000001011000000100000;	//add $s6,$s0,$zero
		17:Instruction<=32'b10001111110010000000000000100000;	//Read2:   lw $t0,8($fp)
		18:Instruction<=32'b00110001000010000000000000001000;	//andi $t0,$t0,8
		19:Instruction<=32'b00010000000010001111111111111101;	//beq $t0,$zero,Read2
		20:Instruction<=32'b10001111110100010000000000011100;	//lw $s1,7($fp)
		21:Instruction<=32'b00000010001000001011100000100000;	//add $s7,$s1,$zero
		22:Instruction<=32'b00000000000000001001000000100000;	//add $s2,$zero,$zero
		23:Instruction<=32'b00000010001100000100000000100010;	//Judge:   sub $t0,$s1,$s0
		24:Instruction<=32'b00010000000010000000000000000110;	//beq $t0,$zero,Result
		25:Instruction<=32'b01001001000000000000000000000011;	//bltz $t0,Minus
		26:Instruction<=32'b00000010000000000100100000100000;	//add $t1,$s0,$zero
		27:Instruction<=32'b00000010001000001000000000100000;	//add $s0,$s1,$zero
		28:Instruction<=32'b00000001001000001000100000100000;	//add $s1,$t1,$zero
		29:Instruction<=32'b00000010000100011000000000100010;	//Minus:   sub $s0,$s0,$s1
		30:Instruction<=32'b00001000000000000000000000010111;	//j Judge
		31:Instruction<=32'b00000000000100011001000000100000;	//Result:   add $s2,$zero,$s1
		32:Instruction<=32'b10101111110100100000000000011000;	//sw $s2,6($fp)
		33:Instruction<=32'b00001000000000000000000000001100;	//j Read1
		34:Instruction<=32'b00100011101111011111111111011100;	//Interrupt:   addi $sp,$sp,-36
		35:Instruction<=32'b10101111101111100000000000100000;	//sw $fp,8($sp)
		36:Instruction<=32'b10101111101101100000000000011100;	//sw $s6,7($sp)
		37:Instruction<=32'b10101111101101110000000000011000;	//sw $s7,6($sp)
		38:Instruction<=32'b10101111101100100000000000010100;	//sw $s2,5($sp)
		39:Instruction<=32'b10101111101110100000000000010000;	//sw $k0,4($sp)
		40:Instruction<=32'b10101111101010000000000000001100;	//sw $t0,3($sp)
		41:Instruction<=32'b10101111101010010000000000001000;	//sw $t1,2($sp)
		42:Instruction<=32'b10101111101100000000000000000100;	//sw $s0,1($sp)
		43:Instruction<=32'b10101111101100010000000000000000;	//sw $s1,0($sp)
		44:Instruction<=32'b10101111110000000000000000001000;	//sw $zero,2($fp)
		45:Instruction<=32'b10001111110010000000000000010100;	//lw $t0,5($fp)
		46:Instruction<=32'b00110001000010010000100000000000;	//andi $t1,$t0,2048
		47:Instruction<=32'b00010000000010010000000000000111;	//beq $t1,$zero,AN2
		48:Instruction<=32'b00110001000010010000010000000000;	//andi $t1,$t0,1024
		49:Instruction<=32'b00010000000010010000000000001000;	//beq $t1,$zero,AN1
		50:Instruction<=32'b00110001000010010000001000000000;	//andi $t1,$t0,512
		51:Instruction<=32'b00010000000010010000000000001001;	//beq $t1,$zero,AN0
		52:Instruction<=32'b00000000000101100100000100000010;	//srl $t0,$s6,4
		53:Instruction<=32'b00100000000010010000011100000000;	//addi $t1,$zero,1792
		54:Instruction<=32'b00001000000000000000000000111111;	//j Trans
		55:Instruction<=32'b00110010110010000000000000001111;	//AN2:   andi $t0,$s6,15
		56:Instruction<=32'b00100000000010010000101100000000;	//addi $t1,$zero,2816
		57:Instruction<=32'b00001000000000000000000000111111;	//j Trans
		58:Instruction<=32'b00000000000101110100000100000010;	//AN1:   srl $t0,$s7,4
		59:Instruction<=32'b00100000000010010000110100000000;	//addi $t1,$zero,3328
		60:Instruction<=32'b00001000000000000000000000111111;	//j Trans
		61:Instruction<=32'b00110010111010000000000000001111;	//AN0:   andi $t0,$s7,15
		62:Instruction<=32'b00100000000010010000111000000000;	//addi $t1,$zero,3584
		63:Instruction<=32'b00010100000010000000000000000010;	//Trans:
		64:Instruction<=32'b00100001001010010000000011000000;	//bne $t0,$zero,One
		65:Instruction<=32'b00001000000000000000000001111011;	//addi $t1,$t1,192
		66:Instruction<=32'b00100001000010001111111111111111;	//j Save
		67:Instruction<=32'b00010100000010000000000000000010;	//One:   addi $t0,$t0,-1
		68:Instruction<=32'b00100001001010010000000011111001;	//bne $t0,$zero,Two
		69:Instruction<=32'b00001000000000000000000001111011;	//addi $t1,$t1,249
		70:Instruction<=32'b00100001000010001111111111111111;	//j Save
		71:Instruction<=32'b00010100000010000000000000000010;	//Two:   addi $t0,$t0,-1
		72:Instruction<=32'b00100001001010010000000010100100;	//bne $t0,$zero,Three
		73:Instruction<=32'b00001000000000000000000001111011;	//addi $t1,$t1,164
		74:Instruction<=32'b00100001000010001111111111111111;	//j Save
		75:Instruction<=32'b00010100000010000000000000000010;	//Three:   addi $t0,$t0,-1
		76:Instruction<=32'b00100001001010010000000010110000;	//bne $t0,$zero,Four
		77:Instruction<=32'b00001000000000000000000001111011;	//addi $t1,$t1,176
		78:Instruction<=32'b00100001000010001111111111111111;	//j Save
		79:Instruction<=32'b00010100000010000000000000000010;	//Four:   addi $t0,$t0,-1
		80:Instruction<=32'b00100001001010010000000010011001;	//bne $t0,$zero,Five
		81:Instruction<=32'b00001000000000000000000001111011;	//addi $t1,$t1,153
		82:Instruction<=32'b00100001000010001111111111111111;	//j Save
		83:Instruction<=32'b00010100000010000000000000000010;	//Five:   addi $t0,$t0,-1
		84:Instruction<=32'b00100001001010010000000010010010;	//bne $t0,$zero,Six
		85:Instruction<=32'b00001000000000000000000001111011;	//addi $t1,$t1,146
		86:Instruction<=32'b00100001000010001111111111111111;	//j Save
		87:Instruction<=32'b00010100000010000000000000000010;	//Six:   addi $t0,$t0,-1
		88:Instruction<=32'b00100001001010010000000010000010;	//bne $t0,$zero,Seven
		89:Instruction<=32'b00001000000000000000000001111011;	//addi $t1,$t1,130
		90:Instruction<=32'b00100001000010001111111111111111;	//j Save
		91:Instruction<=32'b00010100000010000000000000000010;	//Seven:   addi $t0,$t0,-1
		92:Instruction<=32'b00100001001010010000000011111000;	//bne $t0,$zero,Eight
		93:Instruction<=32'b00001000000000000000000001111011;	//addi $t1,$t1,248
		94:Instruction<=32'b00100001000010001111111111111111;	//j Save
		95:Instruction<=32'b00010100000010000000000000000010;	//Eight:   addi $t0,$t0,-1
		96:Instruction<=32'b00100001001010010000000010000000;	//bne $t0,$zero,Nine
		97:Instruction<=32'b00001000000000000000000001111011;	//addi $t1,$t1,128
		98:Instruction<=32'b00100001000010001111111111111111;	//j Save
		99:Instruction<=32'b00010100000010000000000000000010;	//Nine:   addi $t0,$t0,-1
		100:Instruction<=32'b00100001001010010000000010010000;	//bne $t0,$zero,Ten
		101:Instruction<=32'b00001000000000000000000001111011;	//addi $t1,$t1,144
		102:Instruction<=32'b00100001000010001111111111111111;	//j Save
		103:Instruction<=32'b00010100000010000000000000000010;	//Ten:   addi $t0,$t0,-1
		104:Instruction<=32'b00100001001010010000000010001000;	//bne $t0,$zero,Eleven
		105:Instruction<=32'b00001000000000000000000001111011;	//addi $t1,$t1,136
		106:Instruction<=32'b00100001000010001111111111111111;	//j Save
		107:Instruction<=32'b00010100000010000000000000000010;	//Eleven:   addi $t0,$t0,-1
		108:Instruction<=32'b00100001001010010000000010000011;	//bne $t0,$zero,Twelve
		109:Instruction<=32'b00001000000000000000000001111011;	//addi $t1,$t1,131
		110:Instruction<=32'b00100001000010001111111111111111;	//j Save
		111:Instruction<=32'b00010100000010000000000000000010;	//Twelve:   addi $t0,$t0,-1
		112:Instruction<=32'b00100001001010010000000011000110;	//bne $t0,$zero,Thirteen
		113:Instruction<=32'b00001000000000000000000001111011;	//addi $t1,$t1,198
		114:Instruction<=32'b00100001000010001111111111111111;	//j Save
		115:Instruction<=32'b00010100000010000000000000000010;	//Thirteen:   addi $t0,$t0,-1
		116:Instruction<=32'b00100001001010010000000010100001;	//bne $t0,$zero,Fourteen
		117:Instruction<=32'b00001000000000000000000001111011;	//addi $t1,$t1,161
		118:Instruction<=32'b00100001000010001111111111111111;	//j Save
		119:Instruction<=32'b00010100000010000000000000000010;	//Fourteen:   addi $t0,$t0,-1
		120:Instruction<=32'b00100001001010010000000010000110;	//bne $t0,$zero,Fifteen
		121:Instruction<=32'b00001000000000000000000001111011;	//addi $t1,$t1,134
		122:Instruction<=32'b00100001001010010000000010001110;	//j Save
		123:Instruction<=32'b10101111110010010000000000010100;	//Fifteen:   addi $t1,$t1,142
		124:Instruction<=32'b10101111110100100000000000001100;	//Save:   sw $t1,5($fp)
		125:Instruction<=32'b00100000000010000000000000000011;	//sw $s2,3($fp)
		126:Instruction<=32'b10101111110010000000000000001000;	//addi $t0,$zero,3
		127:Instruction<=32'b10001111101100010000000000000000;	//sw $t0,2($fp)
		128:Instruction<=32'b10001111101100000000000000000100;	//lw $s1,0($sp)
		129:Instruction<=32'b10001111101010010000000000001000;	//lw $s0,1($sp)
		130:Instruction<=32'b10001111101010000000000000001100;	//lw $t1,2($sp)
		131:Instruction<=32'b10001111101110100000000000010000;	//lw $t0,3($sp)
		132:Instruction<=32'b10001111101100100000000000010100;	//lw $k0,4($sp)
		133:Instruction<=32'b10001111101101110000000000011000;	//lw $s2,5($sp)
		134:Instruction<=32'b10001111101101100000000000011100;	//lw $s7,6($sp)
		135:Instruction<=32'b10001111101111100000000000100000;	//lw $s6,7($sp)
		136:Instruction<=32'b00100011101111010000000000100100;	//lw $fp,8($sp)
		137:Instruction<=32'b00000011010000000000000000001000;	//addi $sp,$sp,36

		default:Instruction<=32'b00000000000000000000000000000000;
	endcase
endmodule 