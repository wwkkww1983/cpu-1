module Peripheral_S(reset,clk,rd,wr,switch,addr,wdata,rdata,led,digi,IRQ);
input reset;
input clk;
input rd;
input wr;
input [7:0] switch;
input [31:0] addr;
input [31:0] wdata;
output [31:0] rdata;
output [7:0] led;
output [11:0] digi;
output IRQ;

reg [31:0] rdata;
reg [7:0] led;
reg [11:0] digi;
reg [31:0] TH,TL;
reg [2:0] TCON;
assign IRQ=TCON[2];

always@(*) begin
	if(rd) begin
		case(addr)
			32'h40000000: rdata <= TH;			
			32'h40000004: rdata <= TL;			
			32'h40000008: rdata <= {29'b0,TCON};				
			32'h4000000C: rdata <= {24'b0,led};			
			32'h40000010: rdata <= {24'b0,switch};
			32'h40000014: rdata <= {20'b0,digi};
			default: rdata <= 32'b0;
		endcase
	end
	else
		rdata <= 32'b0;
end

always@(posedge reset or posedge clk) begin
	if(reset) begin
		TH <= 32'b0;
		TL <= 32'b0;
		TCON <= 3'b0;
		digi <= 12'b0;	
	end
	else begin
		if(TCON[0]) begin					//timer is enabled
			if(TL==32'hffffffff) begin
				TL <= TH;
				if(TCON[1]) 
					TCON[2] <= 1'b1;		//irq is enabled
			end
			else TL <= TL + 1;
		end
		if(wr) begin
			case(addr)
				32'h40000000: TH <= wdata;
				32'h40000004: TL <= wdata;
				32'h40000008: TCON <= wdata[2:0];		
				32'h4000000C: led <= wdata[7:0];			
				32'h40000014: digi <= wdata[11:0];
				default: ;
			endcase
		end
	end
end
endmodule 